module xillydemo
  (
   input  PCIE_PERST_B_LS,
   input  PCIE_REFCLK_N,
   input  PCIE_REFCLK_P,
   input [7:0] PCIE_RX_N,
   input [7:0] PCIE_RX_P,
   output [3:0] GPIO_LED,
   output [7:0] PCIE_TX_N,
   output [7:0] PCIE_TX_P
   );
   // Clock and quiesce
   wire  bus_clk;
   wire  quiesce;
 
 
   // Wires related to /dev/xillybus_mem_32
   wire  user_r_mem_32_rden;
   wire  user_r_mem_32_empty;
   wire [31:0] user_r_mem_32_data;
   wire  user_r_mem_32_eof;
   wire  user_r_mem_32_open;
   wire  user_w_mem_32_wren;
   wire  user_w_mem_32_full;
   wire [31:0] user_w_mem_32_data;
   wire  user_w_mem_32_open;
   wire [31:0] user_mem_32_addr;
   wire  user_mem_32_addr_update;
 
   // Wires related to /dev/xillybus_read_32
   wire  user_r_read_32_rden;
   wire  user_r_read_32_empty;
   wire [31:0] user_r_read_32_data;
   wire  user_r_read_32_eof;
   wire  user_r_read_32_open;
 
   // Wires related to /dev/xillybus_read_8
   wire  user_r_read_8_rden;
   wire  user_r_read_8_empty;
   wire [7:0] user_r_read_8_data;
   wire  user_r_read_8_eof;
   wire  user_r_read_8_open;
 
   // Wires related to /dev/xillybus_write_32
   wire  user_w_write_32_wren;
   wire  user_w_write_32_full;
   wire [31:0] user_w_write_32_data;
   wire  user_w_write_32_open;
 
   // Wires related to /dev/xillybus_write_8
   wire  user_w_write_8_wren;
   wire  user_w_write_8_full;
   wire [7:0] user_w_write_8_data;
   wire  user_w_write_8_open;
 
 
   xillybus xillybus_ins (
 
     // Ports related to /dev/xillybus_mem_32
     // FPGA to CPU signals:
     .user_r_mem_32_rden(user_r_mem_32_rden),
     .user_r_mem_32_empty(user_r_mem_32_empty),
     .user_r_mem_32_data(user_r_mem_32_data),
     .user_r_mem_32_eof(user_r_mem_32_eof),
     .user_r_mem_32_open(user_r_mem_32_open),
 
     // CPU to FPGA signals:
     .user_w_mem_32_wren(user_w_mem_32_wren),
     .user_w_mem_32_full(user_w_mem_32_full),
     .user_w_mem_32_data(user_w_mem_32_data),
     .user_w_mem_32_open(user_w_mem_32_open),
 
     // Address signals:
     .user_mem_32_addr(user_mem_32_addr),
     .user_mem_32_addr_update(user_mem_32_addr_update),
 
 
     // Ports related to /dev/xillybus_read_32
     // FPGA to CPU signals:
     .user_r_read_32_rden(user_r_read_32_rden),
     .user_r_read_32_empty(user_r_read_32_empty),
     .user_r_read_32_data(user_r_read_32_data),
     .user_r_read_32_eof(user_r_read_32_eof),
     .user_r_read_32_open(user_r_read_32_open),
 
 
     // Ports related to /dev/xillybus_read_8
     // FPGA to CPU signals:
     .user_r_read_8_rden(user_r_read_8_rden),
     .user_r_read_8_empty(user_r_read_8_empty),
     .user_r_read_8_data(user_r_read_8_data),
     .user_r_read_8_eof(user_r_read_8_eof),
     .user_r_read_8_open(user_r_read_8_open),
 
 
     // Ports related to /dev/xillybus_write_32
     // CPU to FPGA signals:
     .user_w_write_32_wren(user_w_write_32_wren),
     .user_w_write_32_full(user_w_write_32_full),
     .user_w_write_32_data(user_w_write_32_data),
     .user_w_write_32_open(user_w_write_32_open),
 
 
     // Ports related to /dev/xillybus_write_8
     // CPU to FPGA signals:
     .user_w_write_8_wren(user_w_write_8_wren),
     .user_w_write_8_full(user_w_write_8_full),
     .user_w_write_8_data(user_w_write_8_data),
     .user_w_write_8_open(user_w_write_8_open),
 
 
     // General signals
     .PCIE_PERST_B_LS(PCIE_PERST_B_LS),
     .PCIE_REFCLK_N(PCIE_REFCLK_N),
     .PCIE_REFCLK_P(PCIE_REFCLK_P),
     .PCIE_RX_N(PCIE_RX_N),
     .PCIE_RX_P(PCIE_RX_P),
     .GPIO_LED(GPIO_LED),
     .PCIE_TX_N(PCIE_TX_N),
     .PCIE_TX_P(PCIE_TX_P),
     .bus_clk(bus_clk),
     .quiesce(quiesce)
   );


   // A simple inferred RAM
   always @(posedge bus_clk)
     begin
	if (user_w_mem_32_wren)
	  demoarray[user_mem_32_addr] <= user_w_mem_32_data;
	
	if (user_r_mem_32_rden)
	  user_r_mem_32_data <= demoarray[user_mem_32_addr];	  
     end

   assign  user_r_mem_32_empty = 0;
   assign  user_r_mem_32_eof = 0;
   assign  user_w_mem_32_full = 0;

   // 32-bit loopback
   fifo_32x512 fifo_32
     (
      .clk(bus_clk),
      .srst(!user_w_write_32_open && !user_r_read_32_open),
      .din(user_w_write_32_data),
      .wr_en(user_w_write_32_wren),
      .rd_en(user_r_read_32_rden),
      .dout(user_r_read_32_data),
      .full(user_w_write_32_full),
      .empty(user_r_read_32_empty)
      );

   assign  user_r_read_32_eof = 0;
   
   // 8-bit loopback
   fifo_8x2048 fifo_8
     (
      .clk(bus_clk),
      .srst(!user_w_write_8_open && !user_r_read_8_open),
      .din(user_w_write_8_data),
      .wr_en(user_w_write_8_wren),
      .rd_en(user_r_read_8_rden),
      .dout(user_r_read_8_data),
      .full(user_w_write_8_full),
      .empty(user_r_read_8_empty)
      );

   assign  user_r_read_8_eof = 0;
   
endmodule
